module ROM_Empate(input [3:0] rom_addr, output [107:0] rom_data);
	always @*
		case (rom_addr)
			0: rom_data = 108'b011111111111111110011111000000111110011111111111111110011111111111111110011111111111111110011111111111111110;
			1: rom_data = 108'b011111111111111110011111100001111110011111111111111110011111111111111110011111111111111110011111111111111110;
			2: rom_data = 108'b011111000000000000011111100001111110011111000000111110011111000000111110000000111111000000011111000000000000;
			3: rom_data = 108'b011111000000000000011111110011111110011111000000111110011111000000111110000000111111000000011111000000000000;
			4: rom_data = 108'b011111000000000000011111110011111110011111000000111110011111000000111110000000111111000000011111000000000000;
			5: rom_data = 108'b011111000000000000011111011110111110011111000000111110011111000000111110000000111111000000011111000000000000;
			6: rom_data = 108'b011111000000000000011111011110111110011111000000111110011111000000111110000000111111000000011111000000000000;
			7: rom_data = 108'b011111111111111000011111011110111110011111111111111110011111111111111110000000111111000000011111111111111000;
			8: rom_data = 108'b011111111111111000011111001100111110011111111111111110011111111111111110000000111111000000011111111111111000;
			9: rom_data = 108'b011111000000000000011111001100111110011111000000000000011111000000111110000000111111000000011111000000000000;
		  10: rom_data = 108'b011111000000000000011111000000111110011111000000000000011111000000111110000000111111000000011111000000000000;
		  11: rom_data = 108'b011111000000000000011111000000111110011111000000000000011111000000111110000000111111000000011111000000000000;
		  12: rom_data = 108'b011111000000000000011111000000111110011111000000000000011111000000111110000000111111000000011111000000000000;
		  13: rom_data = 108'b011111000000000000011111000000111110011111000000000000011111000000111110000000111111000000011111000000000000;
		  14: rom_data = 108'b011111111111111110011111000000111110011111000000000000011111000000111110000000111111000000011111111111111110;
		  15: rom_data = 108'b011111111111111110011111000000111110011111000000000000011111000000111110000000111111000000011111111111111110;

		endcase

endmodule 