module ROM_X_Ganador(input [3:0] rom_addr, output [89:0] rom_data);
	always @*
		case (rom_addr)
			0: rom_data = 90'b011111111111111110011111111111111110011111000000111110011111111111111110011111000000111110;
			1: rom_data = 90'b011111111111111110011111111111111110011111100000111110011111111111111110001111100001111100;
			2: rom_data = 90'b011111000000000000011111111111111110011111110000111110011111000000111110000111110011111000;
			3: rom_data = 90'b011111000000000000011111000000111110011111111000111110011111000000111110000011111111110000;
			4: rom_data = 90'b011111000000000000011111000000111110011111111100111110011111000000111110000001111111100000;
			5: rom_data = 90'b011111000000000000011111000000111110011111111110111110011111000000111110000000111111000000;
			6: rom_data = 90'b011111000000000000011111000000111110011111011111111110011111000000111110000000111111000000;
			7: rom_data = 90'b011111000111111110011111111111111110011111001111111110011111000000111110000001111111100000;
			8: rom_data = 90'b011111000111111110011111111111111110011111000111111110011111000000111110000011111111110000;
			9: rom_data = 90'b011111000111111110011111111111111110011111000011111110011111000000111110000111110011111000;
		  10: rom_data = 90'b011111000000011110011111111111111110011111000001111110011111000000111110001111100001111100;
		  11: rom_data = 90'b011111000000011110011111000000111110011111000000111110011111000000111110011111000000111110;
		  12: rom_data = 90'b011111000000011110011111000000111110011111000000111110011111000000111110011110000000011110;
		  13: rom_data = 90'b011111000000011110011111000000111110011111000000111110011111000000111110011100000000001110;
		  14: rom_data = 90'b011111111111111110011111000000111110011111000000111110011111111111111110011000000000000110;
		  15: rom_data = 90'b011111111111111110011111000000111110011111000000111110011111111111111110010000000000000010;

		endcase

endmodule 