module ROM_Circle_Ganador(input [3:0] rom_addr, output [89:0] rom_data);
	always @*
		case (rom_addr)
			0: rom_data = 90'b011111111111111110011111111111111110011111000000111110011111111111111110000000111111000000;
			1: rom_data = 90'b011111111111111110011111111111111110011111100000111110011111111111111110000011111111110000;
			2: rom_data = 90'b011111000000000000011111111111111110011111110000111110011111000000111110000111111111111000;
			3: rom_data = 90'b011111000000000000011111000000111110011111111000111110011111000000111110001111111111111100;
			4: rom_data = 90'b011111000000000000011111000000111110011111111100111110011111000000111110011111111111111110;
			5: rom_data = 90'b011111000000000000011111000000111110011111111110111110011111000000111110011111111111111110;
			6: rom_data = 90'b011111000000000000011111000000111110011111011111111110011111000000111110011111111111111110;
			7: rom_data = 90'b011111000111111110011111111111111110011111001111111110011111000000111110011111111111111110;
			8: rom_data = 90'b011111000111111110011111111111111110011111000111111110011111000000111110011111111111111110;
			9: rom_data = 90'b011111000111111110011111111111111110011111000011111110011111000000111110011111111111111110;
		  10: rom_data = 90'b011111000000011110011111111111111110011111000001111110011111000000111110011111111111111110;
		  11: rom_data = 90'b011111000000011110011111000000111110011111000000111110011111000000111110011111111111111110;
		  12: rom_data = 90'b011111000000011110011111000000111110011111000000111110011111000000111110001111111111111100;
		  13: rom_data = 90'b011111000000011110011111000000111110011111000000111110011111000000111110000111111111111000;
		  14: rom_data = 90'b011111111111111110011111000000111110011111000000111110011111111111111110000011111111110000;
		  15: rom_data = 90'b011111111111111110011111000000111110011111000000111110011111111111111110000000111111000000;

		endcase

endmodule 