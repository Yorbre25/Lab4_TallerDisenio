//Modulo ROM X
module ROM_X(input [5:0] rom_addr, output [63:0] rom_data);
	always @*
		case (rom_addr)
			0: rom_data = 64'b1111111111111111111100000000000000000000000011111111111111111111;
			1: rom_data = 64'b0111111111111111111110000000000000000000000111111111111111111110;
			2: rom_data = 64'b0011111111111111111111000000000000000000001111111111111111111100;
			3: rom_data = 64'b0001111111111111111111100000000000000000011111111111111111111000;
			4: rom_data = 64'b0000111111111111111111110000000000000000111111111111111111110000;
			5: rom_data = 64'b0000011111111111111111111000000000000001111111111111111111100000;
			6: rom_data = 64'b0000001111111111111111111100000000000011111111111111111111000000;
			7: rom_data = 64'b0000000111111111111111111110000000000111111111111111111110000000;
			8: rom_data = 64'b0000000011111111111111111111000000001111111111111111111100000000;
			9: rom_data = 64'b0000000001111111111111111111100000011111111111111111111000000000;
		  10: rom_data = 64'b0000000000111111111111111111110000111111111111111111110000000000;
		  11: rom_data = 64'b0000000000011111111111111111111001111111111111111111100000000000;
		  12: rom_data = 64'b0000000000001111111111111111111111111111111111111111000000000000;
		  13: rom_data = 64'b0000000000000111111111111111111111111111111111111110000000000000;
		  14: rom_data = 64'b0000000000000011111111111111111111111111111111111100000000000000;
		  15: rom_data = 64'b0000000000000001111111111111111111111111111111111000000000000000;
		  16: rom_data = 64'b0000000000000000111111111111111111111111111111110000000000000000;
		  17: rom_data = 64'b0000000000000000011111111111111111111111111111100000000000000000;
		  18: rom_data = 64'b0000000000000000001111111111111111111111111111000000000000000000;
		  19: rom_data = 64'b0000000000000000000111111111111111111111111110000000000000000000;
		  20: rom_data = 64'b0000000000000000000011111111111111111111111100000000000000000000;
		  21: rom_data = 64'b0000000000000000000001111111111111111111111000000000000000000000;
		  22: rom_data = 64'b0000000000000000000000111111111111111111110000000000000000000000;
		  23: rom_data = 64'b0000000000000000000001111111111111111111111000000000000000000000;
		  24: rom_data = 64'b0000000000000000000011111111111111111111111100000000000000000000;
		  25: rom_data = 64'b0000000000000000000111111111111111111111111110000000000000000000;
		  26: rom_data = 64'b0000000000000000001111111111111111111111111111000000000000000000;
		  27: rom_data = 64'b0000000000000000011111111111111111111111111111100000000000000000;
		  28: rom_data = 64'b0000000000000000111111111111111111111111111111110000000000000000;
		  29: rom_data = 64'b0000000000000001111111111111111111111111111111111000000000000000;
		  30: rom_data = 64'b0000000000000011111111111111111111111111111111111100000000000000;
		  31: rom_data = 64'b0000000000000111111111111111111111111111111111111110000000000000;
		  32: rom_data = 64'b0000000000001111111111111111111111111111111111111111000000000000;
		  33: rom_data = 64'b0000000000011111111111111111111001111111111111111111100000000000;
		  34: rom_data = 64'b0000000000111111111111111111110000111111111111111111110000000000;
		  35: rom_data = 64'b0000000001111111111111111111100000011111111111111111111000000000;
		  36: rom_data = 64'b0000000011111111111111111111000000001111111111111111111100000000;
		  37: rom_data = 64'b0000000111111111111111111110000000000111111111111111111110000000;
		  38: rom_data = 64'b0000001111111111111111111100000000000011111111111111111111000000;
		  39: rom_data = 64'b0000011111111111111111111000000000000001111111111111111111100000;
		  40: rom_data = 64'b0000111111111111111111110000000000000000111111111111111111110000;
		  41: rom_data = 64'b0001111111111111111111100000000000000000011111111111111111111000;
		  42: rom_data = 64'b0011111111111111111111000000000000000000001111111111111111111100;
		  43: rom_data = 64'b0111111111111111111110000000000000000000000111111111111111111110;
		  44: rom_data = 64'b1111111111111111111100000000000000000000000011111111111111111111;
		  45: rom_data = 64'b1111111111111111111000000000000000000000000001111111111111111111;
		  46: rom_data = 64'b1111111111111111110000000000000000000000000000111111111111111111;
		  47: rom_data = 64'b1111111111111111100000000000000000000000000000011111111111111111;
		  48: rom_data = 64'b1111111111111111000000000000000000000000000000001111111111111111;
		  49: rom_data = 64'b1111111111111110000000000000000000000000000000000111111111111111;
		  50: rom_data = 64'b1111111111111100000000000000000000000000000000000011111111111111;
		  51: rom_data = 64'b1111111111111000000000000000000000000000000000000001111111111111;
		  52: rom_data = 64'b1111111111110000000000000000000000000000000000000000111111111111;
		  53: rom_data = 64'b1111111111100000000000000000000000000000000000000000011111111111;
		  54: rom_data = 64'b1111111111000000000000000000000000000000000000000000001111111111;
		  55: rom_data = 64'b1111111110000000000000000000000000000000000000000000000111111111;
		  56: rom_data = 64'b1111111100000000000000000000000000000000000000000000000011111111;
		  57: rom_data = 64'b1111111000000000000000000000000000000000000000000000000001111111;
		  58: rom_data = 64'b1111110000000000000000000000000000000000000000000000000000111111;
		  59: rom_data = 64'b1111100000000000000000000000000000000000000000000000000000011111;
		  60: rom_data = 64'b1111000000000000000000000000000000000000000000000000000000001111;
		  61: rom_data = 64'b1110000000000000000000000000000000000000000000000000000000000111;
		  62: rom_data = 64'b1100000000000000000000000000000000000000000000000000000000000011;
		  63: rom_data = 64'b1000000000000000000000000000000000000000000000000000000000000001;
		  
		endcase

endmodule 