//Probar la FSM de Ganador: Funciona individualmente, pero junto a la matriz no
//Hacer que cuando se gane se reinicie todo el juego
//Reset en matriz no funiciona
//Juntar bien la vara
//Hacer el contador
//La parte random